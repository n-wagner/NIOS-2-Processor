
module NIOSProcessorLab (
	clk_clk);	

	input		clk_clk;
endmodule
