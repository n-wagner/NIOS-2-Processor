
module NIOSProcessor (
	clk_clk);	

	input		clk_clk;
endmodule
